module hehe
fn hoho() {
	println("Hello")
}
