module hehe
pub fn hoho() {
	println("Hello")
}
